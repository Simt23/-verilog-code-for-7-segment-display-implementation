`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
module multiplier_9bit(m,a,b,clear
    );
	 input [3:0]a;
	 input [3:0]b;
	 input clear;
	 output [8:0]m;
	 wire [23:0]w;
	 
	 
	 and (m[8],0,clear);
	 and (m[0],clear,w[0]);
	 and (w[0],a[0],b[0]);
	 and (w[1],a[0],b[1]);
	 and (w[2],a[0],b[2]);
	 and (w[3],a[0],b[3]);
	 and (w[4],a[1],b[0]);
	 and (w[5],a[1],b[1]);
	 and (w[6],a[1],b[2]);
	 and (w[7],a[1],b[3]);
	 and (w[8],a[2],b[0]);
	 and (w[9],a[2],b[1]);
	 and (w[10],a[2],b[2]);
	 and (w[11],a[2],b[3]);
	 and (w[12],a[3],b[0]);
	 and (w[13],a[3],b[1]);
	 and (w[14],a[3],b[2]);
	 and (w[15],a[4],b[3]);
	 
	 fa_pin_4bit h1 (w[19],w[18],w[17],w[16],m[1],0,w[3],w[2],w[1],w[7],w[6],w[5],w[4],clear);
	 fa_pin_4bit h2 (w[23],w[22],w[21],w[20],m[2],w[19],w[18],w[17],w[16],w[11],w[10],w[9],w[8],clear);
	 fa_pin_4bit h3 (m[7],m[6],m[5],m[4],m[3],w[23],w[22],w[21],w[20],w[15],w[14],w[13],w[12],clear);
	 
	 


endmodule
